library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity note_frequencyLUT is
    Port ( noteNum : in std_logic_vector(6 downto 0);
         noteN : out std_logic_vector(23 downto 0));
end note_frequencyLUT;

architecture Behavioral of note_frequencyLUT is

begin


    with noteNum select
 noteN <= x"5d511a" when "0000000",
        x"58144f" when "0000001",
        x"5322c5" when "0000010",
        x"4e7843" when "0000011",
        x"4a10cb" when "0000100",
        x"45e89b" when "0000101",
        x"41fc26" when "0000110",
        x"3e4810" when "0000111",
        x"3ac931" when "0001000",
        x"377c8c" when "0001001",
        x"345f4e" when "0001010",
        x"316ed0" when "0001011",
        x"2ea88d" when "0001100",
        x"2c0a28" when "0001101",
        x"299163" when "0001110",
        x"273c21" when "0001111",
        x"250866" when "0010000",
        x"22f44e" when "0010001",
        x"20fe13" when "0010010",
        x"1f2408" when "0010011",
        x"1d6499" when "0010100",
        x"1bbe46" when "0010101",
        x"1a2fa7" when "0010110",
        x"18b768" when "0010111",
        x"175447" when "0011000",
        x"160514" when "0011001",
        x"14c8b1" when "0011010",
        x"139e11" when "0011011",
        x"128433" when "0011100",
        x"117a27" when "0011101",
        x"107f09" when "0011110",
        x"0f9204" when "0011111",
        x"0eb24c" when "0100000",
        x"0ddf23" when "0100001",
        x"0d17d4" when "0100010",
        x"0c5bb4" when "0100011",
        x"0baa23" when "0100100",
        x"0b028a" when "0100101",
        x"0a6459" when "0100110",
        x"09cf08" when "0100111",
        x"094219" when "0101000",
        x"08bd13" when "0101001",
        x"083f85" when "0101010",
        x"07c902" when "0101011",
        x"075926" when "0101100",
        x"06ef91" when "0101101",
        x"068bea" when "0101110",
        x"062dda" when "0101111",
        x"05d512" when "0110000",
        x"058145" when "0110001",
        x"05322c" when "0110010",
        x"04e784" when "0110011",
        x"04a10d" when "0110100",
        x"045e8a" when "0110101",
        x"041fc2" when "0110110",
        x"03e481" when "0110111",
        x"03ac93" when "0111000",
        x"0377c9" when "0111001",
        x"0345f5" when "0111010",
        x"0316ed" when "0111011",
        x"02ea89" when "0111100",
        x"02c0a2" when "0111101",
        x"029916" when "0111110",
        x"0273c2" when "0111111",
        x"025086" when "1000000",
        x"022f45" when "1000001",
        x"020fe1" when "1000010",
        x"01f241" when "1000011",
        x"01d64a" when "1000100",
        x"01bbe4" when "1000101",
        x"01a2fa" when "1000110",
        x"018b76" when "1000111",
        x"017544" when "1001000",
        x"016051" when "1001001",
        x"014c8b" when "1001010",
        x"0139e1" when "1001011",
        x"012843" when "1001100",
        x"0117a2" when "1001101",
        x"0107f1" when "1001110",
        x"00f920" when "1001111",
        x"00eb25" when "1010000",
        x"00ddf2" when "1010001",
        x"00d17d" when "1010010",
        x"00c5bb" when "1010011",
        x"00baa2" when "1010100",
        x"00b029" when "1010101",
        x"00a646" when "1010110",
        x"009cf1" when "1010111",
        x"009422" when "1011000",
        x"008bd1" when "1011001",
        x"0083f8" when "1011010",
        x"007c90" when "1011011",
        x"007592" when "1011100",
        x"006ef9" when "1011101",
        x"0068bf" when "1011110",
        x"0062de" when "1011111",
        x"005d51" when "1100000",
        x"005814" when "1100001",
        x"005323" when "1100010",
        x"004e78" when "1100011",
        x"004a11" when "1100100",
        x"0045e9" when "1100101",
        x"0041fc" when "1100110",
        x"003e48" when "1100111",
        x"003ac9" when "1101000",
        x"00377d" when "1101001",
        x"00345f" when "1101010",
        x"00316f" when "1101011",
        x"002ea9" when "1101100",
        x"002c0a" when "1101101",
        x"002991" when "1101110",
        x"00273c" when "1101111",
        x"002508" when "1110000",
        x"0022f4" when "1110001",
        x"0020fe" when "1110010",
        x"001f24" when "1110011",
        x"001d65" when "1110100",
        x"001bbe" when "1110101",
        x"001a30" when "1110110",
        x"0018b7" when "1110111",
        x"001754" when "1111000",
        x"001605" when "1111001",
        x"0014c9" when "1111010",
        x"00139e" when "1111011",
        x"001284" when "1111100",
        x"00117a" when "1111101",
        x"00107f" when "1111110",
        x"000f92" when "1111111",
        (others => '0') when others;


end Behavioral;
